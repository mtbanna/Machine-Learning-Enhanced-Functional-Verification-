package tests_package;
     `include "bus_request_test.sv"
     `include "basic_transfer_single_master_single_slave_test.sv"
     `include "default_master_and_slave_test.sv"
     `include "basic_read_single_master_single_slave_test.sv"
     `include "reset_assertion_and_deassertion_test.sv"
     `include "arbitration_and_hold_idle_state_test.sv"
     `include "locked_write_single_master_single_slave_test.sv"
endpackage 