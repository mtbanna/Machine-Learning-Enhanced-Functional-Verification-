package coverages_package;
     `include "bus_request_coverage.sv"
     `include "basic_transfer_single_master_single_slave_coverage.sv"
     `include "default_master_and_slave_coverage.sv"
     `include "basic_read_single_master_single_slave_coverage.sv"
     `include "reset_assertion_and_deassertion_coverage.sv"
     `include "arbitration_and_hold_idle_state_coverage.sv"
     `include "locked_write_single_master_single_slave_coverage.sv"
endpackage 