package sequences_package;
     `include "bus_request_sequence.sv"
     `include "basic_transfer_single_master_single_slave_sequence.sv"
     `include "default_master_and_slave_sequence.sv"
     `include "basic_read_single_master_single_slave_sequence.sv"
     `include "reset_assertion_and_deassertion_sequence.sv"
     `include "arbitration_and_hold_idle_state_sequence.sv"
     `include "locked_write_single_master_single_slave_sequence.sv"
endpackage 