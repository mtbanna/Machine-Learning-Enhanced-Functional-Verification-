package scoreboards_package;
     `include "bus_request_scoreboard.sv"
     `include "basic_transfer_single_master_single_slave_scoreboard.sv"
     `include "default_master_and_slave_scoreboard.sv"
     `include "basic_read_single_master_single_slave_scoreboard.sv"
     `include "reset_assertion_and_deassertion_scoreboard.sv"
     `include "arbitration_and_hold_idle_state_scoreboard.sv"
     `include "locked_write_single_master_single_slave_scoreboard.sv"     
endpackage 